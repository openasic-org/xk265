//--------------------------------------------------------------------
//
//  Filename    : ime_ver_mem.v
//  Author      : Huang Leilei
//  Created     : 2018-06-18
//  Description : vertical memory in ime module
//
//--------------------------------------------------------------------
`include "enc_defines.v"
module ime_ver_mem(
  // global
  clk             ,
  rstn            ,
  // cfg_i
  rotate_i        ,
  downsample_i    ,
  // wr_if
  wr_dir_i        ,
  wr_ena_i        ,
  wr_adr_x_i      ,
  wr_adr_y_i      ,
  wr_dat_i        ,
  // rd_if
  rd_ena_i        ,
  rd_adr_x_i      ,
  rd_adr_y_i      ,
  rd_dat_o
  );


//*** PARAMETER ****************************************************************


//*** INPUT/OUTPUT *************************************************************

  // global
  input                                      clk              ;
  input                                      rstn             ;
  // ctrl_if
  input                                      rotate_i         ;
  input                                      downsample_i     ;
  // ref_rd
  input      [2                    -1 :0]    wr_dir_i         ;
  input      [1                    -1 :0]    wr_ena_i         ;
  input      [`IME_MV_WIDTH_Y         :0]    wr_adr_x_i       ;
  input      [`IME_MV_WIDTH_X         :0]    wr_adr_y_i       ;
  input      [`IME_PIXEL_WIDTH*1024-1 :0]    wr_dat_i         ;
  // ref_wr
  input                                      rd_ena_i         ;
  input      [`IME_MV_WIDTH_Y         :0]    rd_adr_x_i       ;
  input      [`IME_MV_WIDTH_X         :0]    rd_adr_y_i       ;
  output reg [`IME_PIXEL_WIDTH*32  -1 :0]    rd_dat_o         ;


//*** REG/WIRE ***************************************************************

  // rotater
  reg        [2                    -1 :0]    rot_cnt_r        ;
  wire                                       rot_done_w       ;

  // write
  reg        [`IME_PIXEL_WIDTH*128 -1 :0]    wr_ena_w         ;
  reg        [`IME_MV_WIDTH_X         :0]    wr_adr_w         ;
  reg        [`IME_PIXEL_WIDTH*128 -1 :0]    wr_dat_w         ;
  wire       [`IME_PIXEL_WIDTH*32  -1 :0]    wr_dat_hor_w     ;
  wire       [`IME_PIXEL_WIDTH*32  -1 :0]    wr_dat_ver_w     ;

  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_00_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_01_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_02_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_03_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_04_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_05_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_06_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_07_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_08_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_09_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_10_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_11_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_12_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_13_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_14_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_15_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_16_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_17_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_18_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_19_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_20_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_21_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_22_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_23_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_24_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_25_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_26_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_27_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_28_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_29_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_30_31_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_00_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_01_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_02_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_03_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_04_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_05_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_06_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_07_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_08_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_09_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_10_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_11_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_12_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_13_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_14_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_15_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_16_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_17_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_18_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_19_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_20_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_21_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_22_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_23_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_24_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_25_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_26_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_27_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_28_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_29_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_30_w   ;
  wire       [`IME_PIXEL_WIDTH     -1 :0]    wr_dat_31_31_w   ;

  // read
  reg        [`IME_MV_WIDTH_X         :0]    rd_adr_w         ;
  wire       [`IME_PIXEL_WIDTH*128 -1 :0]    rd_dat_w         ;
  wire       [`IME_PIXEL_WIDTH*128 -1 :0]    rd_dat_shif_w    ;

  reg        [`IME_MV_WIDTH_Y         :0]    rd_adr_x         ;

  // adr
  wire       [`IME_MV_WIDTH_X         :0]    adr_w            ;


//*** MAIN BODY ****************************************************************

//--- GLOBAL ---------------------------
  // rotater
  always @(posedge clk or negedge rstn ) begin
    if( !rstn ) begin
      rot_cnt_r <= 0 ;
    end
    else begin
      if( rotate_i ) begin
        if( rot_done_w ) begin
          rot_cnt_r <= 0 ;
        end
        else begin
          rot_cnt_r <= rot_cnt_r + 1 ;
        end
      end
    end
  end

  assign rot_done_w = rot_cnt_r == 2 ;


//--- WRITE ----------------------------
  // wr_ena_w
  always @(*) begin
           wr_ena_w = 0    ;
    if ( wr_ena_i ) begin
      case( wr_adr_x_i[6:5] )
        0  : wr_ena_w = { {(`IME_PIXEL_WIDTH*32){1'b1}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} };
        1  : wr_ena_w = { {(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b1}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} };
        2  : wr_ena_w = { {(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b1}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} };
        3  : wr_ena_w = { {(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b0}} ,{(`IME_PIXEL_WIDTH*32){1'b1}} };
      endcase
    end
    else begin
      wr_ena_w = 0 ;
    end
  end

  // wr_adr_w
  always @(*) begin
                         wr_adr_w = 0 ;
    case( rot_cnt_r )
      0 : begin          wr_adr_w = wr_adr_y_i ;
      end
      1 : begin    case( wr_adr_y_i[7:5] )
                     0 : wr_adr_w = { 3'd2 ,wr_adr_y_i[4:0] };
                     1 : wr_adr_w = { 3'd3 ,wr_adr_y_i[4:0] };
                     2 : wr_adr_w = { 3'd4 ,wr_adr_y_i[4:0] };
                     3 : wr_adr_w = { 3'd5 ,wr_adr_y_i[4:0] };
                     4 : wr_adr_w = { 3'd0 ,wr_adr_y_i[4:0] };
                     5 : wr_adr_w = { 3'd1 ,wr_adr_y_i[4:0] };
                   endcase
      end
      2 : begin    case( wr_adr_y_i[7:5] )
                     0 : wr_adr_w = { 3'd4 ,wr_adr_y_i[4:0] };
                     1 : wr_adr_w = { 3'd5 ,wr_adr_y_i[4:0] };
                     2 : wr_adr_w = { 3'd0 ,wr_adr_y_i[4:0] };
                     3 : wr_adr_w = { 3'd1 ,wr_adr_y_i[4:0] };
                     4 : wr_adr_w = { 3'd2 ,wr_adr_y_i[4:0] };
                     5 : wr_adr_w = { 3'd3 ,wr_adr_y_i[4:0] };
                   endcase
      end
    endcase
  end

  // wr_dat_w
  always @(*) begin
                       wr_dat_w = {{(`IME_PIXEL_WIDTH*128){1'b0}}} ;
    case( wr_dir_i )
      `IME_DIR_DOWN  : wr_dat_w = {{4{wr_dat_hor_w}}} ;
      `IME_DIR_RIGHT : wr_dat_w = {{4{wr_dat_ver_w}}} ;
    endcase
  end

  // wr_dat_hor_w    
  assign wr_dat_hor_w = { wr_dat_00_00_w,wr_dat_00_01_w,wr_dat_00_02_w,wr_dat_00_03_w,wr_dat_00_04_w,wr_dat_00_05_w,wr_dat_00_06_w,wr_dat_00_07_w,wr_dat_00_08_w,wr_dat_00_09_w,wr_dat_00_10_w,wr_dat_00_11_w,wr_dat_00_12_w,wr_dat_00_13_w,wr_dat_00_14_w,wr_dat_00_15_w,wr_dat_00_16_w,wr_dat_00_17_w,wr_dat_00_18_w,wr_dat_00_19_w,wr_dat_00_20_w,wr_dat_00_21_w,wr_dat_00_22_w,wr_dat_00_23_w,wr_dat_00_24_w,wr_dat_00_25_w,wr_dat_00_26_w,wr_dat_00_27_w,wr_dat_00_28_w,wr_dat_00_29_w,wr_dat_00_30_w,wr_dat_00_31_w };

  // wr_dat_ver_w    
  assign wr_dat_ver_w = { wr_dat_00_00_w,wr_dat_01_00_w,wr_dat_02_00_w,wr_dat_03_00_w,wr_dat_04_00_w,wr_dat_05_00_w,wr_dat_06_00_w,wr_dat_07_00_w,wr_dat_08_00_w,wr_dat_09_00_w,wr_dat_10_00_w,wr_dat_11_00_w,wr_dat_12_00_w,wr_dat_13_00_w,wr_dat_14_00_w,wr_dat_15_00_w,wr_dat_16_00_w,wr_dat_17_00_w,wr_dat_18_00_w,wr_dat_19_00_w,wr_dat_20_00_w,wr_dat_21_00_w,wr_dat_22_00_w,wr_dat_23_00_w,wr_dat_24_00_w,wr_dat_25_00_w,wr_dat_26_00_w,wr_dat_27_00_w,wr_dat_28_00_w,wr_dat_29_00_w,wr_dat_30_00_w,wr_dat_31_00_w };

  // wr_dat_xx_xx_w
  assign { wr_dat_00_00_w
          ,wr_dat_00_01_w
          ,wr_dat_00_02_w
          ,wr_dat_00_03_w
          ,wr_dat_00_04_w
          ,wr_dat_00_05_w
          ,wr_dat_00_06_w
          ,wr_dat_00_07_w
          ,wr_dat_00_08_w
          ,wr_dat_00_09_w
          ,wr_dat_00_10_w
          ,wr_dat_00_11_w
          ,wr_dat_00_12_w
          ,wr_dat_00_13_w
          ,wr_dat_00_14_w
          ,wr_dat_00_15_w
          ,wr_dat_00_16_w
          ,wr_dat_00_17_w
          ,wr_dat_00_18_w
          ,wr_dat_00_19_w
          ,wr_dat_00_20_w
          ,wr_dat_00_21_w
          ,wr_dat_00_22_w
          ,wr_dat_00_23_w
          ,wr_dat_00_24_w
          ,wr_dat_00_25_w
          ,wr_dat_00_26_w
          ,wr_dat_00_27_w
          ,wr_dat_00_28_w
          ,wr_dat_00_29_w
          ,wr_dat_00_30_w
          ,wr_dat_00_31_w
          ,wr_dat_01_00_w
          ,wr_dat_01_01_w
          ,wr_dat_01_02_w
          ,wr_dat_01_03_w
          ,wr_dat_01_04_w
          ,wr_dat_01_05_w
          ,wr_dat_01_06_w
          ,wr_dat_01_07_w
          ,wr_dat_01_08_w
          ,wr_dat_01_09_w
          ,wr_dat_01_10_w
          ,wr_dat_01_11_w
          ,wr_dat_01_12_w
          ,wr_dat_01_13_w
          ,wr_dat_01_14_w
          ,wr_dat_01_15_w
          ,wr_dat_01_16_w
          ,wr_dat_01_17_w
          ,wr_dat_01_18_w
          ,wr_dat_01_19_w
          ,wr_dat_01_20_w
          ,wr_dat_01_21_w
          ,wr_dat_01_22_w
          ,wr_dat_01_23_w
          ,wr_dat_01_24_w
          ,wr_dat_01_25_w
          ,wr_dat_01_26_w
          ,wr_dat_01_27_w
          ,wr_dat_01_28_w
          ,wr_dat_01_29_w
          ,wr_dat_01_30_w
          ,wr_dat_01_31_w
          ,wr_dat_02_00_w
          ,wr_dat_02_01_w
          ,wr_dat_02_02_w
          ,wr_dat_02_03_w
          ,wr_dat_02_04_w
          ,wr_dat_02_05_w
          ,wr_dat_02_06_w
          ,wr_dat_02_07_w
          ,wr_dat_02_08_w
          ,wr_dat_02_09_w
          ,wr_dat_02_10_w
          ,wr_dat_02_11_w
          ,wr_dat_02_12_w
          ,wr_dat_02_13_w
          ,wr_dat_02_14_w
          ,wr_dat_02_15_w
          ,wr_dat_02_16_w
          ,wr_dat_02_17_w
          ,wr_dat_02_18_w
          ,wr_dat_02_19_w
          ,wr_dat_02_20_w
          ,wr_dat_02_21_w
          ,wr_dat_02_22_w
          ,wr_dat_02_23_w
          ,wr_dat_02_24_w
          ,wr_dat_02_25_w
          ,wr_dat_02_26_w
          ,wr_dat_02_27_w
          ,wr_dat_02_28_w
          ,wr_dat_02_29_w
          ,wr_dat_02_30_w
          ,wr_dat_02_31_w
          ,wr_dat_03_00_w
          ,wr_dat_03_01_w
          ,wr_dat_03_02_w
          ,wr_dat_03_03_w
          ,wr_dat_03_04_w
          ,wr_dat_03_05_w
          ,wr_dat_03_06_w
          ,wr_dat_03_07_w
          ,wr_dat_03_08_w
          ,wr_dat_03_09_w
          ,wr_dat_03_10_w
          ,wr_dat_03_11_w
          ,wr_dat_03_12_w
          ,wr_dat_03_13_w
          ,wr_dat_03_14_w
          ,wr_dat_03_15_w
          ,wr_dat_03_16_w
          ,wr_dat_03_17_w
          ,wr_dat_03_18_w
          ,wr_dat_03_19_w
          ,wr_dat_03_20_w
          ,wr_dat_03_21_w
          ,wr_dat_03_22_w
          ,wr_dat_03_23_w
          ,wr_dat_03_24_w
          ,wr_dat_03_25_w
          ,wr_dat_03_26_w
          ,wr_dat_03_27_w
          ,wr_dat_03_28_w
          ,wr_dat_03_29_w
          ,wr_dat_03_30_w
          ,wr_dat_03_31_w
          ,wr_dat_04_00_w
          ,wr_dat_04_01_w
          ,wr_dat_04_02_w
          ,wr_dat_04_03_w
          ,wr_dat_04_04_w
          ,wr_dat_04_05_w
          ,wr_dat_04_06_w
          ,wr_dat_04_07_w
          ,wr_dat_04_08_w
          ,wr_dat_04_09_w
          ,wr_dat_04_10_w
          ,wr_dat_04_11_w
          ,wr_dat_04_12_w
          ,wr_dat_04_13_w
          ,wr_dat_04_14_w
          ,wr_dat_04_15_w
          ,wr_dat_04_16_w
          ,wr_dat_04_17_w
          ,wr_dat_04_18_w
          ,wr_dat_04_19_w
          ,wr_dat_04_20_w
          ,wr_dat_04_21_w
          ,wr_dat_04_22_w
          ,wr_dat_04_23_w
          ,wr_dat_04_24_w
          ,wr_dat_04_25_w
          ,wr_dat_04_26_w
          ,wr_dat_04_27_w
          ,wr_dat_04_28_w
          ,wr_dat_04_29_w
          ,wr_dat_04_30_w
          ,wr_dat_04_31_w
          ,wr_dat_05_00_w
          ,wr_dat_05_01_w
          ,wr_dat_05_02_w
          ,wr_dat_05_03_w
          ,wr_dat_05_04_w
          ,wr_dat_05_05_w
          ,wr_dat_05_06_w
          ,wr_dat_05_07_w
          ,wr_dat_05_08_w
          ,wr_dat_05_09_w
          ,wr_dat_05_10_w
          ,wr_dat_05_11_w
          ,wr_dat_05_12_w
          ,wr_dat_05_13_w
          ,wr_dat_05_14_w
          ,wr_dat_05_15_w
          ,wr_dat_05_16_w
          ,wr_dat_05_17_w
          ,wr_dat_05_18_w
          ,wr_dat_05_19_w
          ,wr_dat_05_20_w
          ,wr_dat_05_21_w
          ,wr_dat_05_22_w
          ,wr_dat_05_23_w
          ,wr_dat_05_24_w
          ,wr_dat_05_25_w
          ,wr_dat_05_26_w
          ,wr_dat_05_27_w
          ,wr_dat_05_28_w
          ,wr_dat_05_29_w
          ,wr_dat_05_30_w
          ,wr_dat_05_31_w
          ,wr_dat_06_00_w
          ,wr_dat_06_01_w
          ,wr_dat_06_02_w
          ,wr_dat_06_03_w
          ,wr_dat_06_04_w
          ,wr_dat_06_05_w
          ,wr_dat_06_06_w
          ,wr_dat_06_07_w
          ,wr_dat_06_08_w
          ,wr_dat_06_09_w
          ,wr_dat_06_10_w
          ,wr_dat_06_11_w
          ,wr_dat_06_12_w
          ,wr_dat_06_13_w
          ,wr_dat_06_14_w
          ,wr_dat_06_15_w
          ,wr_dat_06_16_w
          ,wr_dat_06_17_w
          ,wr_dat_06_18_w
          ,wr_dat_06_19_w
          ,wr_dat_06_20_w
          ,wr_dat_06_21_w
          ,wr_dat_06_22_w
          ,wr_dat_06_23_w
          ,wr_dat_06_24_w
          ,wr_dat_06_25_w
          ,wr_dat_06_26_w
          ,wr_dat_06_27_w
          ,wr_dat_06_28_w
          ,wr_dat_06_29_w
          ,wr_dat_06_30_w
          ,wr_dat_06_31_w
          ,wr_dat_07_00_w
          ,wr_dat_07_01_w
          ,wr_dat_07_02_w
          ,wr_dat_07_03_w
          ,wr_dat_07_04_w
          ,wr_dat_07_05_w
          ,wr_dat_07_06_w
          ,wr_dat_07_07_w
          ,wr_dat_07_08_w
          ,wr_dat_07_09_w
          ,wr_dat_07_10_w
          ,wr_dat_07_11_w
          ,wr_dat_07_12_w
          ,wr_dat_07_13_w
          ,wr_dat_07_14_w
          ,wr_dat_07_15_w
          ,wr_dat_07_16_w
          ,wr_dat_07_17_w
          ,wr_dat_07_18_w
          ,wr_dat_07_19_w
          ,wr_dat_07_20_w
          ,wr_dat_07_21_w
          ,wr_dat_07_22_w
          ,wr_dat_07_23_w
          ,wr_dat_07_24_w
          ,wr_dat_07_25_w
          ,wr_dat_07_26_w
          ,wr_dat_07_27_w
          ,wr_dat_07_28_w
          ,wr_dat_07_29_w
          ,wr_dat_07_30_w
          ,wr_dat_07_31_w
          ,wr_dat_08_00_w
          ,wr_dat_08_01_w
          ,wr_dat_08_02_w
          ,wr_dat_08_03_w
          ,wr_dat_08_04_w
          ,wr_dat_08_05_w
          ,wr_dat_08_06_w
          ,wr_dat_08_07_w
          ,wr_dat_08_08_w
          ,wr_dat_08_09_w
          ,wr_dat_08_10_w
          ,wr_dat_08_11_w
          ,wr_dat_08_12_w
          ,wr_dat_08_13_w
          ,wr_dat_08_14_w
          ,wr_dat_08_15_w
          ,wr_dat_08_16_w
          ,wr_dat_08_17_w
          ,wr_dat_08_18_w
          ,wr_dat_08_19_w
          ,wr_dat_08_20_w
          ,wr_dat_08_21_w
          ,wr_dat_08_22_w
          ,wr_dat_08_23_w
          ,wr_dat_08_24_w
          ,wr_dat_08_25_w
          ,wr_dat_08_26_w
          ,wr_dat_08_27_w
          ,wr_dat_08_28_w
          ,wr_dat_08_29_w
          ,wr_dat_08_30_w
          ,wr_dat_08_31_w
          ,wr_dat_09_00_w
          ,wr_dat_09_01_w
          ,wr_dat_09_02_w
          ,wr_dat_09_03_w
          ,wr_dat_09_04_w
          ,wr_dat_09_05_w
          ,wr_dat_09_06_w
          ,wr_dat_09_07_w
          ,wr_dat_09_08_w
          ,wr_dat_09_09_w
          ,wr_dat_09_10_w
          ,wr_dat_09_11_w
          ,wr_dat_09_12_w
          ,wr_dat_09_13_w
          ,wr_dat_09_14_w
          ,wr_dat_09_15_w
          ,wr_dat_09_16_w
          ,wr_dat_09_17_w
          ,wr_dat_09_18_w
          ,wr_dat_09_19_w
          ,wr_dat_09_20_w
          ,wr_dat_09_21_w
          ,wr_dat_09_22_w
          ,wr_dat_09_23_w
          ,wr_dat_09_24_w
          ,wr_dat_09_25_w
          ,wr_dat_09_26_w
          ,wr_dat_09_27_w
          ,wr_dat_09_28_w
          ,wr_dat_09_29_w
          ,wr_dat_09_30_w
          ,wr_dat_09_31_w
          ,wr_dat_10_00_w
          ,wr_dat_10_01_w
          ,wr_dat_10_02_w
          ,wr_dat_10_03_w
          ,wr_dat_10_04_w
          ,wr_dat_10_05_w
          ,wr_dat_10_06_w
          ,wr_dat_10_07_w
          ,wr_dat_10_08_w
          ,wr_dat_10_09_w
          ,wr_dat_10_10_w
          ,wr_dat_10_11_w
          ,wr_dat_10_12_w
          ,wr_dat_10_13_w
          ,wr_dat_10_14_w
          ,wr_dat_10_15_w
          ,wr_dat_10_16_w
          ,wr_dat_10_17_w
          ,wr_dat_10_18_w
          ,wr_dat_10_19_w
          ,wr_dat_10_20_w
          ,wr_dat_10_21_w
          ,wr_dat_10_22_w
          ,wr_dat_10_23_w
          ,wr_dat_10_24_w
          ,wr_dat_10_25_w
          ,wr_dat_10_26_w
          ,wr_dat_10_27_w
          ,wr_dat_10_28_w
          ,wr_dat_10_29_w
          ,wr_dat_10_30_w
          ,wr_dat_10_31_w
          ,wr_dat_11_00_w
          ,wr_dat_11_01_w
          ,wr_dat_11_02_w
          ,wr_dat_11_03_w
          ,wr_dat_11_04_w
          ,wr_dat_11_05_w
          ,wr_dat_11_06_w
          ,wr_dat_11_07_w
          ,wr_dat_11_08_w
          ,wr_dat_11_09_w
          ,wr_dat_11_10_w
          ,wr_dat_11_11_w
          ,wr_dat_11_12_w
          ,wr_dat_11_13_w
          ,wr_dat_11_14_w
          ,wr_dat_11_15_w
          ,wr_dat_11_16_w
          ,wr_dat_11_17_w
          ,wr_dat_11_18_w
          ,wr_dat_11_19_w
          ,wr_dat_11_20_w
          ,wr_dat_11_21_w
          ,wr_dat_11_22_w
          ,wr_dat_11_23_w
          ,wr_dat_11_24_w
          ,wr_dat_11_25_w
          ,wr_dat_11_26_w
          ,wr_dat_11_27_w
          ,wr_dat_11_28_w
          ,wr_dat_11_29_w
          ,wr_dat_11_30_w
          ,wr_dat_11_31_w
          ,wr_dat_12_00_w
          ,wr_dat_12_01_w
          ,wr_dat_12_02_w
          ,wr_dat_12_03_w
          ,wr_dat_12_04_w
          ,wr_dat_12_05_w
          ,wr_dat_12_06_w
          ,wr_dat_12_07_w
          ,wr_dat_12_08_w
          ,wr_dat_12_09_w
          ,wr_dat_12_10_w
          ,wr_dat_12_11_w
          ,wr_dat_12_12_w
          ,wr_dat_12_13_w
          ,wr_dat_12_14_w
          ,wr_dat_12_15_w
          ,wr_dat_12_16_w
          ,wr_dat_12_17_w
          ,wr_dat_12_18_w
          ,wr_dat_12_19_w
          ,wr_dat_12_20_w
          ,wr_dat_12_21_w
          ,wr_dat_12_22_w
          ,wr_dat_12_23_w
          ,wr_dat_12_24_w
          ,wr_dat_12_25_w
          ,wr_dat_12_26_w
          ,wr_dat_12_27_w
          ,wr_dat_12_28_w
          ,wr_dat_12_29_w
          ,wr_dat_12_30_w
          ,wr_dat_12_31_w
          ,wr_dat_13_00_w
          ,wr_dat_13_01_w
          ,wr_dat_13_02_w
          ,wr_dat_13_03_w
          ,wr_dat_13_04_w
          ,wr_dat_13_05_w
          ,wr_dat_13_06_w
          ,wr_dat_13_07_w
          ,wr_dat_13_08_w
          ,wr_dat_13_09_w
          ,wr_dat_13_10_w
          ,wr_dat_13_11_w
          ,wr_dat_13_12_w
          ,wr_dat_13_13_w
          ,wr_dat_13_14_w
          ,wr_dat_13_15_w
          ,wr_dat_13_16_w
          ,wr_dat_13_17_w
          ,wr_dat_13_18_w
          ,wr_dat_13_19_w
          ,wr_dat_13_20_w
          ,wr_dat_13_21_w
          ,wr_dat_13_22_w
          ,wr_dat_13_23_w
          ,wr_dat_13_24_w
          ,wr_dat_13_25_w
          ,wr_dat_13_26_w
          ,wr_dat_13_27_w
          ,wr_dat_13_28_w
          ,wr_dat_13_29_w
          ,wr_dat_13_30_w
          ,wr_dat_13_31_w
          ,wr_dat_14_00_w
          ,wr_dat_14_01_w
          ,wr_dat_14_02_w
          ,wr_dat_14_03_w
          ,wr_dat_14_04_w
          ,wr_dat_14_05_w
          ,wr_dat_14_06_w
          ,wr_dat_14_07_w
          ,wr_dat_14_08_w
          ,wr_dat_14_09_w
          ,wr_dat_14_10_w
          ,wr_dat_14_11_w
          ,wr_dat_14_12_w
          ,wr_dat_14_13_w
          ,wr_dat_14_14_w
          ,wr_dat_14_15_w
          ,wr_dat_14_16_w
          ,wr_dat_14_17_w
          ,wr_dat_14_18_w
          ,wr_dat_14_19_w
          ,wr_dat_14_20_w
          ,wr_dat_14_21_w
          ,wr_dat_14_22_w
          ,wr_dat_14_23_w
          ,wr_dat_14_24_w
          ,wr_dat_14_25_w
          ,wr_dat_14_26_w
          ,wr_dat_14_27_w
          ,wr_dat_14_28_w
          ,wr_dat_14_29_w
          ,wr_dat_14_30_w
          ,wr_dat_14_31_w
          ,wr_dat_15_00_w
          ,wr_dat_15_01_w
          ,wr_dat_15_02_w
          ,wr_dat_15_03_w
          ,wr_dat_15_04_w
          ,wr_dat_15_05_w
          ,wr_dat_15_06_w
          ,wr_dat_15_07_w
          ,wr_dat_15_08_w
          ,wr_dat_15_09_w
          ,wr_dat_15_10_w
          ,wr_dat_15_11_w
          ,wr_dat_15_12_w
          ,wr_dat_15_13_w
          ,wr_dat_15_14_w
          ,wr_dat_15_15_w
          ,wr_dat_15_16_w
          ,wr_dat_15_17_w
          ,wr_dat_15_18_w
          ,wr_dat_15_19_w
          ,wr_dat_15_20_w
          ,wr_dat_15_21_w
          ,wr_dat_15_22_w
          ,wr_dat_15_23_w
          ,wr_dat_15_24_w
          ,wr_dat_15_25_w
          ,wr_dat_15_26_w
          ,wr_dat_15_27_w
          ,wr_dat_15_28_w
          ,wr_dat_15_29_w
          ,wr_dat_15_30_w
          ,wr_dat_15_31_w
          ,wr_dat_16_00_w
          ,wr_dat_16_01_w
          ,wr_dat_16_02_w
          ,wr_dat_16_03_w
          ,wr_dat_16_04_w
          ,wr_dat_16_05_w
          ,wr_dat_16_06_w
          ,wr_dat_16_07_w
          ,wr_dat_16_08_w
          ,wr_dat_16_09_w
          ,wr_dat_16_10_w
          ,wr_dat_16_11_w
          ,wr_dat_16_12_w
          ,wr_dat_16_13_w
          ,wr_dat_16_14_w
          ,wr_dat_16_15_w
          ,wr_dat_16_16_w
          ,wr_dat_16_17_w
          ,wr_dat_16_18_w
          ,wr_dat_16_19_w
          ,wr_dat_16_20_w
          ,wr_dat_16_21_w
          ,wr_dat_16_22_w
          ,wr_dat_16_23_w
          ,wr_dat_16_24_w
          ,wr_dat_16_25_w
          ,wr_dat_16_26_w
          ,wr_dat_16_27_w
          ,wr_dat_16_28_w
          ,wr_dat_16_29_w
          ,wr_dat_16_30_w
          ,wr_dat_16_31_w
          ,wr_dat_17_00_w
          ,wr_dat_17_01_w
          ,wr_dat_17_02_w
          ,wr_dat_17_03_w
          ,wr_dat_17_04_w
          ,wr_dat_17_05_w
          ,wr_dat_17_06_w
          ,wr_dat_17_07_w
          ,wr_dat_17_08_w
          ,wr_dat_17_09_w
          ,wr_dat_17_10_w
          ,wr_dat_17_11_w
          ,wr_dat_17_12_w
          ,wr_dat_17_13_w
          ,wr_dat_17_14_w
          ,wr_dat_17_15_w
          ,wr_dat_17_16_w
          ,wr_dat_17_17_w
          ,wr_dat_17_18_w
          ,wr_dat_17_19_w
          ,wr_dat_17_20_w
          ,wr_dat_17_21_w
          ,wr_dat_17_22_w
          ,wr_dat_17_23_w
          ,wr_dat_17_24_w
          ,wr_dat_17_25_w
          ,wr_dat_17_26_w
          ,wr_dat_17_27_w
          ,wr_dat_17_28_w
          ,wr_dat_17_29_w
          ,wr_dat_17_30_w
          ,wr_dat_17_31_w
          ,wr_dat_18_00_w
          ,wr_dat_18_01_w
          ,wr_dat_18_02_w
          ,wr_dat_18_03_w
          ,wr_dat_18_04_w
          ,wr_dat_18_05_w
          ,wr_dat_18_06_w
          ,wr_dat_18_07_w
          ,wr_dat_18_08_w
          ,wr_dat_18_09_w
          ,wr_dat_18_10_w
          ,wr_dat_18_11_w
          ,wr_dat_18_12_w
          ,wr_dat_18_13_w
          ,wr_dat_18_14_w
          ,wr_dat_18_15_w
          ,wr_dat_18_16_w
          ,wr_dat_18_17_w
          ,wr_dat_18_18_w
          ,wr_dat_18_19_w
          ,wr_dat_18_20_w
          ,wr_dat_18_21_w
          ,wr_dat_18_22_w
          ,wr_dat_18_23_w
          ,wr_dat_18_24_w
          ,wr_dat_18_25_w
          ,wr_dat_18_26_w
          ,wr_dat_18_27_w
          ,wr_dat_18_28_w
          ,wr_dat_18_29_w
          ,wr_dat_18_30_w
          ,wr_dat_18_31_w
          ,wr_dat_19_00_w
          ,wr_dat_19_01_w
          ,wr_dat_19_02_w
          ,wr_dat_19_03_w
          ,wr_dat_19_04_w
          ,wr_dat_19_05_w
          ,wr_dat_19_06_w
          ,wr_dat_19_07_w
          ,wr_dat_19_08_w
          ,wr_dat_19_09_w
          ,wr_dat_19_10_w
          ,wr_dat_19_11_w
          ,wr_dat_19_12_w
          ,wr_dat_19_13_w
          ,wr_dat_19_14_w
          ,wr_dat_19_15_w
          ,wr_dat_19_16_w
          ,wr_dat_19_17_w
          ,wr_dat_19_18_w
          ,wr_dat_19_19_w
          ,wr_dat_19_20_w
          ,wr_dat_19_21_w
          ,wr_dat_19_22_w
          ,wr_dat_19_23_w
          ,wr_dat_19_24_w
          ,wr_dat_19_25_w
          ,wr_dat_19_26_w
          ,wr_dat_19_27_w
          ,wr_dat_19_28_w
          ,wr_dat_19_29_w
          ,wr_dat_19_30_w
          ,wr_dat_19_31_w
          ,wr_dat_20_00_w
          ,wr_dat_20_01_w
          ,wr_dat_20_02_w
          ,wr_dat_20_03_w
          ,wr_dat_20_04_w
          ,wr_dat_20_05_w
          ,wr_dat_20_06_w
          ,wr_dat_20_07_w
          ,wr_dat_20_08_w
          ,wr_dat_20_09_w
          ,wr_dat_20_10_w
          ,wr_dat_20_11_w
          ,wr_dat_20_12_w
          ,wr_dat_20_13_w
          ,wr_dat_20_14_w
          ,wr_dat_20_15_w
          ,wr_dat_20_16_w
          ,wr_dat_20_17_w
          ,wr_dat_20_18_w
          ,wr_dat_20_19_w
          ,wr_dat_20_20_w
          ,wr_dat_20_21_w
          ,wr_dat_20_22_w
          ,wr_dat_20_23_w
          ,wr_dat_20_24_w
          ,wr_dat_20_25_w
          ,wr_dat_20_26_w
          ,wr_dat_20_27_w
          ,wr_dat_20_28_w
          ,wr_dat_20_29_w
          ,wr_dat_20_30_w
          ,wr_dat_20_31_w
          ,wr_dat_21_00_w
          ,wr_dat_21_01_w
          ,wr_dat_21_02_w
          ,wr_dat_21_03_w
          ,wr_dat_21_04_w
          ,wr_dat_21_05_w
          ,wr_dat_21_06_w
          ,wr_dat_21_07_w
          ,wr_dat_21_08_w
          ,wr_dat_21_09_w
          ,wr_dat_21_10_w
          ,wr_dat_21_11_w
          ,wr_dat_21_12_w
          ,wr_dat_21_13_w
          ,wr_dat_21_14_w
          ,wr_dat_21_15_w
          ,wr_dat_21_16_w
          ,wr_dat_21_17_w
          ,wr_dat_21_18_w
          ,wr_dat_21_19_w
          ,wr_dat_21_20_w
          ,wr_dat_21_21_w
          ,wr_dat_21_22_w
          ,wr_dat_21_23_w
          ,wr_dat_21_24_w
          ,wr_dat_21_25_w
          ,wr_dat_21_26_w
          ,wr_dat_21_27_w
          ,wr_dat_21_28_w
          ,wr_dat_21_29_w
          ,wr_dat_21_30_w
          ,wr_dat_21_31_w
          ,wr_dat_22_00_w
          ,wr_dat_22_01_w
          ,wr_dat_22_02_w
          ,wr_dat_22_03_w
          ,wr_dat_22_04_w
          ,wr_dat_22_05_w
          ,wr_dat_22_06_w
          ,wr_dat_22_07_w
          ,wr_dat_22_08_w
          ,wr_dat_22_09_w
          ,wr_dat_22_10_w
          ,wr_dat_22_11_w
          ,wr_dat_22_12_w
          ,wr_dat_22_13_w
          ,wr_dat_22_14_w
          ,wr_dat_22_15_w
          ,wr_dat_22_16_w
          ,wr_dat_22_17_w
          ,wr_dat_22_18_w
          ,wr_dat_22_19_w
          ,wr_dat_22_20_w
          ,wr_dat_22_21_w
          ,wr_dat_22_22_w
          ,wr_dat_22_23_w
          ,wr_dat_22_24_w
          ,wr_dat_22_25_w
          ,wr_dat_22_26_w
          ,wr_dat_22_27_w
          ,wr_dat_22_28_w
          ,wr_dat_22_29_w
          ,wr_dat_22_30_w
          ,wr_dat_22_31_w
          ,wr_dat_23_00_w
          ,wr_dat_23_01_w
          ,wr_dat_23_02_w
          ,wr_dat_23_03_w
          ,wr_dat_23_04_w
          ,wr_dat_23_05_w
          ,wr_dat_23_06_w
          ,wr_dat_23_07_w
          ,wr_dat_23_08_w
          ,wr_dat_23_09_w
          ,wr_dat_23_10_w
          ,wr_dat_23_11_w
          ,wr_dat_23_12_w
          ,wr_dat_23_13_w
          ,wr_dat_23_14_w
          ,wr_dat_23_15_w
          ,wr_dat_23_16_w
          ,wr_dat_23_17_w
          ,wr_dat_23_18_w
          ,wr_dat_23_19_w
          ,wr_dat_23_20_w
          ,wr_dat_23_21_w
          ,wr_dat_23_22_w
          ,wr_dat_23_23_w
          ,wr_dat_23_24_w
          ,wr_dat_23_25_w
          ,wr_dat_23_26_w
          ,wr_dat_23_27_w
          ,wr_dat_23_28_w
          ,wr_dat_23_29_w
          ,wr_dat_23_30_w
          ,wr_dat_23_31_w
          ,wr_dat_24_00_w
          ,wr_dat_24_01_w
          ,wr_dat_24_02_w
          ,wr_dat_24_03_w
          ,wr_dat_24_04_w
          ,wr_dat_24_05_w
          ,wr_dat_24_06_w
          ,wr_dat_24_07_w
          ,wr_dat_24_08_w
          ,wr_dat_24_09_w
          ,wr_dat_24_10_w
          ,wr_dat_24_11_w
          ,wr_dat_24_12_w
          ,wr_dat_24_13_w
          ,wr_dat_24_14_w
          ,wr_dat_24_15_w
          ,wr_dat_24_16_w
          ,wr_dat_24_17_w
          ,wr_dat_24_18_w
          ,wr_dat_24_19_w
          ,wr_dat_24_20_w
          ,wr_dat_24_21_w
          ,wr_dat_24_22_w
          ,wr_dat_24_23_w
          ,wr_dat_24_24_w
          ,wr_dat_24_25_w
          ,wr_dat_24_26_w
          ,wr_dat_24_27_w
          ,wr_dat_24_28_w
          ,wr_dat_24_29_w
          ,wr_dat_24_30_w
          ,wr_dat_24_31_w
          ,wr_dat_25_00_w
          ,wr_dat_25_01_w
          ,wr_dat_25_02_w
          ,wr_dat_25_03_w
          ,wr_dat_25_04_w
          ,wr_dat_25_05_w
          ,wr_dat_25_06_w
          ,wr_dat_25_07_w
          ,wr_dat_25_08_w
          ,wr_dat_25_09_w
          ,wr_dat_25_10_w
          ,wr_dat_25_11_w
          ,wr_dat_25_12_w
          ,wr_dat_25_13_w
          ,wr_dat_25_14_w
          ,wr_dat_25_15_w
          ,wr_dat_25_16_w
          ,wr_dat_25_17_w
          ,wr_dat_25_18_w
          ,wr_dat_25_19_w
          ,wr_dat_25_20_w
          ,wr_dat_25_21_w
          ,wr_dat_25_22_w
          ,wr_dat_25_23_w
          ,wr_dat_25_24_w
          ,wr_dat_25_25_w
          ,wr_dat_25_26_w
          ,wr_dat_25_27_w
          ,wr_dat_25_28_w
          ,wr_dat_25_29_w
          ,wr_dat_25_30_w
          ,wr_dat_25_31_w
          ,wr_dat_26_00_w
          ,wr_dat_26_01_w
          ,wr_dat_26_02_w
          ,wr_dat_26_03_w
          ,wr_dat_26_04_w
          ,wr_dat_26_05_w
          ,wr_dat_26_06_w
          ,wr_dat_26_07_w
          ,wr_dat_26_08_w
          ,wr_dat_26_09_w
          ,wr_dat_26_10_w
          ,wr_dat_26_11_w
          ,wr_dat_26_12_w
          ,wr_dat_26_13_w
          ,wr_dat_26_14_w
          ,wr_dat_26_15_w
          ,wr_dat_26_16_w
          ,wr_dat_26_17_w
          ,wr_dat_26_18_w
          ,wr_dat_26_19_w
          ,wr_dat_26_20_w
          ,wr_dat_26_21_w
          ,wr_dat_26_22_w
          ,wr_dat_26_23_w
          ,wr_dat_26_24_w
          ,wr_dat_26_25_w
          ,wr_dat_26_26_w
          ,wr_dat_26_27_w
          ,wr_dat_26_28_w
          ,wr_dat_26_29_w
          ,wr_dat_26_30_w
          ,wr_dat_26_31_w
          ,wr_dat_27_00_w
          ,wr_dat_27_01_w
          ,wr_dat_27_02_w
          ,wr_dat_27_03_w
          ,wr_dat_27_04_w
          ,wr_dat_27_05_w
          ,wr_dat_27_06_w
          ,wr_dat_27_07_w
          ,wr_dat_27_08_w
          ,wr_dat_27_09_w
          ,wr_dat_27_10_w
          ,wr_dat_27_11_w
          ,wr_dat_27_12_w
          ,wr_dat_27_13_w
          ,wr_dat_27_14_w
          ,wr_dat_27_15_w
          ,wr_dat_27_16_w
          ,wr_dat_27_17_w
          ,wr_dat_27_18_w
          ,wr_dat_27_19_w
          ,wr_dat_27_20_w
          ,wr_dat_27_21_w
          ,wr_dat_27_22_w
          ,wr_dat_27_23_w
          ,wr_dat_27_24_w
          ,wr_dat_27_25_w
          ,wr_dat_27_26_w
          ,wr_dat_27_27_w
          ,wr_dat_27_28_w
          ,wr_dat_27_29_w
          ,wr_dat_27_30_w
          ,wr_dat_27_31_w
          ,wr_dat_28_00_w
          ,wr_dat_28_01_w
          ,wr_dat_28_02_w
          ,wr_dat_28_03_w
          ,wr_dat_28_04_w
          ,wr_dat_28_05_w
          ,wr_dat_28_06_w
          ,wr_dat_28_07_w
          ,wr_dat_28_08_w
          ,wr_dat_28_09_w
          ,wr_dat_28_10_w
          ,wr_dat_28_11_w
          ,wr_dat_28_12_w
          ,wr_dat_28_13_w
          ,wr_dat_28_14_w
          ,wr_dat_28_15_w
          ,wr_dat_28_16_w
          ,wr_dat_28_17_w
          ,wr_dat_28_18_w
          ,wr_dat_28_19_w
          ,wr_dat_28_20_w
          ,wr_dat_28_21_w
          ,wr_dat_28_22_w
          ,wr_dat_28_23_w
          ,wr_dat_28_24_w
          ,wr_dat_28_25_w
          ,wr_dat_28_26_w
          ,wr_dat_28_27_w
          ,wr_dat_28_28_w
          ,wr_dat_28_29_w
          ,wr_dat_28_30_w
          ,wr_dat_28_31_w
          ,wr_dat_29_00_w
          ,wr_dat_29_01_w
          ,wr_dat_29_02_w
          ,wr_dat_29_03_w
          ,wr_dat_29_04_w
          ,wr_dat_29_05_w
          ,wr_dat_29_06_w
          ,wr_dat_29_07_w
          ,wr_dat_29_08_w
          ,wr_dat_29_09_w
          ,wr_dat_29_10_w
          ,wr_dat_29_11_w
          ,wr_dat_29_12_w
          ,wr_dat_29_13_w
          ,wr_dat_29_14_w
          ,wr_dat_29_15_w
          ,wr_dat_29_16_w
          ,wr_dat_29_17_w
          ,wr_dat_29_18_w
          ,wr_dat_29_19_w
          ,wr_dat_29_20_w
          ,wr_dat_29_21_w
          ,wr_dat_29_22_w
          ,wr_dat_29_23_w
          ,wr_dat_29_24_w
          ,wr_dat_29_25_w
          ,wr_dat_29_26_w
          ,wr_dat_29_27_w
          ,wr_dat_29_28_w
          ,wr_dat_29_29_w
          ,wr_dat_29_30_w
          ,wr_dat_29_31_w
          ,wr_dat_30_00_w
          ,wr_dat_30_01_w
          ,wr_dat_30_02_w
          ,wr_dat_30_03_w
          ,wr_dat_30_04_w
          ,wr_dat_30_05_w
          ,wr_dat_30_06_w
          ,wr_dat_30_07_w
          ,wr_dat_30_08_w
          ,wr_dat_30_09_w
          ,wr_dat_30_10_w
          ,wr_dat_30_11_w
          ,wr_dat_30_12_w
          ,wr_dat_30_13_w
          ,wr_dat_30_14_w
          ,wr_dat_30_15_w
          ,wr_dat_30_16_w
          ,wr_dat_30_17_w
          ,wr_dat_30_18_w
          ,wr_dat_30_19_w
          ,wr_dat_30_20_w
          ,wr_dat_30_21_w
          ,wr_dat_30_22_w
          ,wr_dat_30_23_w
          ,wr_dat_30_24_w
          ,wr_dat_30_25_w
          ,wr_dat_30_26_w
          ,wr_dat_30_27_w
          ,wr_dat_30_28_w
          ,wr_dat_30_29_w
          ,wr_dat_30_30_w
          ,wr_dat_30_31_w
          ,wr_dat_31_00_w
          ,wr_dat_31_01_w
          ,wr_dat_31_02_w
          ,wr_dat_31_03_w
          ,wr_dat_31_04_w
          ,wr_dat_31_05_w
          ,wr_dat_31_06_w
          ,wr_dat_31_07_w
          ,wr_dat_31_08_w
          ,wr_dat_31_09_w
          ,wr_dat_31_10_w
          ,wr_dat_31_11_w
          ,wr_dat_31_12_w
          ,wr_dat_31_13_w
          ,wr_dat_31_14_w
          ,wr_dat_31_15_w
          ,wr_dat_31_16_w
          ,wr_dat_31_17_w
          ,wr_dat_31_18_w
          ,wr_dat_31_19_w
          ,wr_dat_31_20_w
          ,wr_dat_31_21_w
          ,wr_dat_31_22_w
          ,wr_dat_31_23_w
          ,wr_dat_31_24_w
          ,wr_dat_31_25_w
          ,wr_dat_31_26_w
          ,wr_dat_31_27_w
          ,wr_dat_31_28_w
          ,wr_dat_31_29_w
          ,wr_dat_31_30_w
          ,wr_dat_31_31_w
         } = wr_dat_i ;


//--- READ -----------------------------
  // rd_adr_w
  always @(*) begin
                         rd_adr_w = 0 ;
    case( rot_cnt_r )
      0 : begin          rd_adr_w = rd_adr_y_i ;
      end
      1 : begin    case( rd_adr_y_i[7:5] )
                     0 : rd_adr_w = { 3'd2 ,rd_adr_y_i[4:0] };
                     1 : rd_adr_w = { 3'd3 ,rd_adr_y_i[4:0] };
                     2 : rd_adr_w = { 3'd4 ,rd_adr_y_i[4:0] };
                     3 : rd_adr_w = { 3'd5 ,rd_adr_y_i[4:0] };
                     4 : rd_adr_w = { 3'd0 ,rd_adr_y_i[4:0] };
                     5 : rd_adr_w = { 3'd1 ,rd_adr_y_i[4:0] };
                   endcase
      end
      2 : begin    case( rd_adr_y_i[7:5] )
                     0 : rd_adr_w = { 3'd4 ,rd_adr_y_i[4:0] };
                     1 : rd_adr_w = { 3'd5 ,rd_adr_y_i[4:0] };
                     2 : rd_adr_w = { 3'd0 ,rd_adr_y_i[4:0] };
                     3 : rd_adr_w = { 3'd1 ,rd_adr_y_i[4:0] };
                     4 : rd_adr_w = { 3'd2 ,rd_adr_y_i[4:0] };
                     5 : rd_adr_w = { 3'd3 ,rd_adr_y_i[4:0] };
                   endcase
      end
    endcase
  end


//--- MEMORY ---------------------------
  // adr
  assign adr_w = wr_ena_i ? wr_adr_w : rd_adr_w ;

  // inst
  ram_sp_be_192x512 vertical_memory(
    // global
    .clk         ( clk         ),
    // address
    .adr_i       ( adr_w       ),
    // write
    .wr_ena_i    ( wr_ena_w    ),
    .wr_dat_i    ( wr_dat_w    ),
    // read
    .rd_ena_i    ( rd_ena_i    ),
    .rd_dat_o    ( rd_dat_w    )
    );

  // rd_dat_o
  always @ (posedge clk or negedge rstn) begin
    if (~rstn) begin
      rd_adr_x <= 'd0;
    end
    else begin
      rd_adr_x <= rd_adr_x_i;
    end
  end

  assign rd_dat_shif_w = rd_dat_w << ( rd_adr_x*`IME_PIXEL_WIDTH ) ; 
  
  always @(posedge clk or negedge rstn ) begin
    if( !rstn ) begin
      rd_dat_o <= 0 ;
    end
    else begin
      if (downsample_i)
        rd_dat_o <= { rd_dat_shif_w[`IME_PIXEL_WIDTH*128-1:`IME_PIXEL_WIDTH*127],rd_dat_shif_w[`IME_PIXEL_WIDTH*126-1:`IME_PIXEL_WIDTH*125],rd_dat_shif_w[`IME_PIXEL_WIDTH*124-1:`IME_PIXEL_WIDTH*123],rd_dat_shif_w[`IME_PIXEL_WIDTH*122-1:`IME_PIXEL_WIDTH*121],rd_dat_shif_w[`IME_PIXEL_WIDTH*120-1:`IME_PIXEL_WIDTH*119],
                      rd_dat_shif_w[`IME_PIXEL_WIDTH*118-1:`IME_PIXEL_WIDTH*117],rd_dat_shif_w[`IME_PIXEL_WIDTH*116-1:`IME_PIXEL_WIDTH*115],rd_dat_shif_w[`IME_PIXEL_WIDTH*114-1:`IME_PIXEL_WIDTH*113],rd_dat_shif_w[`IME_PIXEL_WIDTH*112-1:`IME_PIXEL_WIDTH*111],rd_dat_shif_w[`IME_PIXEL_WIDTH*110-1:`IME_PIXEL_WIDTH*109],
                      rd_dat_shif_w[`IME_PIXEL_WIDTH*108-1:`IME_PIXEL_WIDTH*107],rd_dat_shif_w[`IME_PIXEL_WIDTH*106-1:`IME_PIXEL_WIDTH*105],rd_dat_shif_w[`IME_PIXEL_WIDTH*104-1:`IME_PIXEL_WIDTH*103],rd_dat_shif_w[`IME_PIXEL_WIDTH*102-1:`IME_PIXEL_WIDTH*101],rd_dat_shif_w[`IME_PIXEL_WIDTH*100-1:`IME_PIXEL_WIDTH* 99],
                      rd_dat_shif_w[`IME_PIXEL_WIDTH* 98-1:`IME_PIXEL_WIDTH* 97],rd_dat_shif_w[`IME_PIXEL_WIDTH* 96-1:`IME_PIXEL_WIDTH* 95],rd_dat_shif_w[`IME_PIXEL_WIDTH* 94-1:`IME_PIXEL_WIDTH* 93],rd_dat_shif_w[`IME_PIXEL_WIDTH* 92-1:`IME_PIXEL_WIDTH* 91],rd_dat_shif_w[`IME_PIXEL_WIDTH* 90-1:`IME_PIXEL_WIDTH* 89],
                      rd_dat_shif_w[`IME_PIXEL_WIDTH* 88-1:`IME_PIXEL_WIDTH* 87],rd_dat_shif_w[`IME_PIXEL_WIDTH* 86-1:`IME_PIXEL_WIDTH* 85],rd_dat_shif_w[`IME_PIXEL_WIDTH* 84-1:`IME_PIXEL_WIDTH* 83],rd_dat_shif_w[`IME_PIXEL_WIDTH* 82-1:`IME_PIXEL_WIDTH* 81],rd_dat_shif_w[`IME_PIXEL_WIDTH* 80-1:`IME_PIXEL_WIDTH* 79],
                      rd_dat_shif_w[`IME_PIXEL_WIDTH* 78-1:`IME_PIXEL_WIDTH* 77],rd_dat_shif_w[`IME_PIXEL_WIDTH* 76-1:`IME_PIXEL_WIDTH* 75],rd_dat_shif_w[`IME_PIXEL_WIDTH* 74-1:`IME_PIXEL_WIDTH* 73],rd_dat_shif_w[`IME_PIXEL_WIDTH* 72-1:`IME_PIXEL_WIDTH* 71],rd_dat_shif_w[`IME_PIXEL_WIDTH* 70-1:`IME_PIXEL_WIDTH* 69],
                      rd_dat_shif_w[`IME_PIXEL_WIDTH* 68-1:`IME_PIXEL_WIDTH* 67],rd_dat_shif_w[`IME_PIXEL_WIDTH* 66-1:`IME_PIXEL_WIDTH* 65] } ;
      else
        rd_dat_o <=   rd_dat_shif_w[`IME_PIXEL_WIDTH*128-1:`IME_PIXEL_WIDTH*96] ; 
    end
  end

endmodule
